// -*-C++-*-
// Purpose: CDL file to generate netCDF test file 
// Usage:
// ncgen -k netCDF-4 -b -o test_01.nc test_01.cdl

netcdf test_01 {
 dimensions:
  latitude=2;
  longitude=4;
  level=3;
  time=unlimited; 
  dimension_latitude=2;
  dimension_longitude=4;
  dimension_level=3;
  dim_time=unlimited;
 variables:
  double time(time);
  float latitude(latitude);
  float longitude(longitude);
  float level(level);  
  float scl;
  int one_dmn_var_crd(time);
  int one_dmn_var(dim_time);
  float two_dmn_var_crd(latitude,longitude);
  float two_dmn_var(dimension_latitude,dimension_longitude);
  float three_dmn_var_crd(level,latitude,longitude);
  float three_dmn_var(dimension_level,dimension_latitude,dimension_longitude);
 data:
  latitude=-90,90;
  longitude=15,25,35,45;
  level=1000,2000,3000;
  time=10,20,30,40,50,60,70,80,90,100;
  scl=1.0;
  one_dmn_var_crd=1,2,3,4,5,6,7,8,9,10; 
  one_dmn_var=1,2,3,4,5,6,7,8,9,10; 
  two_dmn_var_crd=1,2,3,4,5,6,7,8;
  two_dmn_var=1,2,3,4,5,6,7,8;
  three_dmn_var_crd=1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24;
  three_dmn_var=1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24;
}
