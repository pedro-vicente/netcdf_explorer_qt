// -*-C++-*-
// Purpose: CDL file to generate netCDF test file 
// Usage:
// ncgen -k netCDF-4 -b -o test_02.nc test_02.cdl

netcdf test_02 {
 dimensions:
  time=2;
  level=3; //layers
  latitude=4; //rows
  longitude=5; //columns
 variables:
  float time(time);
  float level(level);
  float latitude(latitude);
  float longitude(longitude);
  float four_dmn_var_crd(time,level,latitude,longitude);
 data:
  time=1,2;
  level=1000,2000,3000;
  latitude=10,20,30,40;
  longitude=100,200,300,400,500;
  four_dmn_var_crd=1, 2, 3, 4, 5, 6, 7, 8, 9, 10,11,12,13,14,15,16,17,18,19,20, // time 0, level 0
                   21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40, // time 0, level 1
                   41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60, // time 0, level 2
                   61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80, // time 1, level 0
                   81,82,83,84,85,86,87,88,99,90,91,92,93,94,95,96,97,98,99,100, // time 2, level 1
                   101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120; // time 3, level 2
 
   
}
