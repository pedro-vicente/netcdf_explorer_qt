// -*-C++-*-
// Purpose: CDL file to generate netCDF test file 
// Usage:
// ncgen -k netCDF-4 -b -o test_03.nc test_03.cdl

netcdf test_02 {
 dimensions:
  gravity=2;
  time=3;
  level=4; //layers
  latitude=2; //rows
  longitude=3; //columns
 variables:
  float gravity(gravity);
  float time(time);
  float level(level);
  float latitude(latitude);
  float longitude(longitude);
  float five_dmn_var_crd(gravity,time,level,latitude,longitude);
 data:
  gravity=1,2;
  time=10,20,30;
  level=1000,2000,3000,4000;
  latitude=100,200;
  longitude=100,200,300;
  five_dmn_var_crd=1, 2, 3, 4, 5, 6,  
                   7, 8, 9, 10,11,12, 
                   13,14,15,16,17,18, 
                   19,20,21,22,23,24, 
                   25,26,27,28,29,30, 
                   31,32,33,34,35,36, 
                   37,38,39,40,41,42, 
                   43,44,45,46,47,48,
                   49,50,51,52,53,54,
                   55,56,57,58,59,60,
                   61,62,63,64,65,66,
                   67,68,69,70,71,72,
                   73,74,75,76,77,78,
                   79,80,81,82,83,84,
                   85,86,87,88,89,90,
                   91,92,93,94,95,96,
                   97,98,99,100,101,102,
                   103,104,105,106,107,108,
                   109,110,111,112,113,114,
                   115,116,117,118,119,120,
                   121,122,123,124,125,126,
                   127,128,129,130,131,132,
                   133,134,135,136,137,138,
                   139,140,141,142,143,144; 
}
